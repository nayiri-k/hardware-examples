module test;
  reg clock = 1;
  reg reset = 1;
  reg[0:0] clock = 0;
  wire[0:0] clock_delay;
  assign  clock_delay = clock;
  reg[0:0] reset = 0;
  wire[0:0] reset_delay;
  assign  reset_delay = reset;
  reg[0:0] io_load = 0;
  wire[0:0] io_load_delay;
  assign  io_load_delay = io_load;
  reg[15:0] io_b = 0;
  wire[15:0] io_b_delay;
  assign  io_b_delay = io_b;
  reg[15:0] io_a = 0;
  wire[15:0] io_a_delay;
  assign  io_a_delay = io_a;
  wire[0:0] io_valid_delay;
  wire[0:0] io_valid;
  assign  io_valid = io_valid_delay;
  wire[15:0] io_out_delay;
  wire[15:0] io_out;
  assign  io_out = io_out_delay;
  always #`CLOCK_PERIOD clock = ~clock;
  reg vcdon = 0;
  reg [1023:0] vcdfile = 0;
  reg [1023:0] vpdfile = 0;

  /*** DUT instantiation ***/
  GCD GCD(
    .clock(clock),
    .reset(reset),
    .clock(clock_delay),
    .reset(reset_delay),
    .io_load(io_load_delay),
    .io_b(io_b_delay),
    .io_a(io_a_delay),
    .io_valid(io_valid_delay),
    .io_out(io_out_delay)  );

  initial begin
    $init_rsts(reset);
    $init_ins(clock, reset, io_load, io_b, io_a);
    $init_outs(io_valid, io_out);
    $init_sigs(GCD);
    /*** VCD & VPD dump ***/
    if ($value$plusargs("vcdfile=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, GCD);
      $dumpoff;
      vcdon = 0;
    end
    if ($value$plusargs("waveform=%s", vpdfile)) begin
      $vcdplusfile(vpdfile);
    end else begin
      $vcdplusfile("generated-src/basic/GCD/GCD.vpd");
    end
    if ($test$plusargs("vpdmem")) begin
      $vcdplusmemon;
    end
    $vcdpluson(0);
  end

  always @(negedge clock) begin
    if (vcdfile && reset) begin
      $dumpoff;
      vcdon = 0;
    end
    else if (vcdfile && !vcdon) begin
      $dumpon;
      vcdon = 1;
    end
     $tick();
    $vcdplusflush;
  end

endmodule
